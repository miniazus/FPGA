//////////////////////////////////////////////////////////////////////////////////
// Company/Author: Viet Ha Nguyen
// Module Name   : UnbiasedRounding
// Date          : November 10, 2025
// Description   : Performs unbiased rounding (round-half-to-even) for fixed-point
//                 numbers. The module truncates the lower bits of the input, applies
//                 rounding based on the truncated portion, and saturates the output
//                 if rounding causes overflow. Supports both signed and unsigned
//                 inputs, and handles fractional or integer rounding modes.
//
// Parameters:
//   DATA_WIDTH_IN_MAX  : Width of the input number
//   DATA_WIDTH_OUT : Width of the output number
//   IS_SIGNED      : Set to 1 for signed input/output, 0 for unsigned
//
// Inputs:
//   clk  : Clock signal for synchronous output
//   ena  : Enable signal to update output
//  din_t  : Input number of DATA_WIDTH_IN_MAX bits
//
// Outputs:
//   dout : Rounded and saturated output of DATA_WIDTH_OUT bits
//
// Features:
//   - Unbiased rounding (round-half-to-even) for tie cases
//   - Saturation to prevent overflow on output
//   - Synthesizable for FPGA/ASIC
//   - Pass-through mode when output width equals input width
//
// Using:
// UnbiasedRounding #(.WIDTH_IN_MAX(...),.WIDTH_OUT(...),.IS_SIGNED(...))
//                 (.clk(...),.ena(...),.width_in(...),.din(...),.dout(...));
//
//////////////////////////////////////////////////////////////////////////////////

module UnbiasedRounding_v2 #(
    parameter int  WIDTH_IN_MAX = 19,
    parameter int  WIDTH_OUT    = 16,
    parameter bit  IS_SIGNED    = 1      // 0 = unsigned, 1 = signed
)
(
    input  logic clk, ena,
    input  logic [7:0] width_in,
    input  logic [WIDTH_IN_MAX-1 :0] din,
    output logic [WIDTH_OUT-1:0]     dout
);
    // Difference in width between input and output
    localparam int                         DIFFWIDTH   = WIDTH_IN_MAX-WIDTH_OUT;
    // Maximum and minimum output values for saturation
    localparam signed   [WIDTH_OUT-1:0]    MAXVALunsigned = {(WIDTH_OUT){1'b1}};
    localparam signed   [WIDTH_OUT-1:0]    MAXVALsigned   = {1'b0, {(WIDTH_OUT-1){1'b1}}};
    localparam signed   [WIDTH_OUT-1:0]    MINVALsigned   = {1'b1, {(WIDTH_OUT-1){1'b0}}};
    // Halfway value used for round-half-to-even
    localparam unsigned [DIFFWIDTH-1:0]    FRAC05      = 1 << (DIFFWIDTH-1);


    logic [WIDTH_IN_MAX-1 :0] din_t;

    generate
        if (IS_SIGNED)
            assign din_t = din <<< (WIDTH_IN_MAX - width_in);
        else
            assign din_t = din <<  (WIDTH_IN_MAX - width_in);
    endgenerate


    generate
        // Check parameter validity
        if (WIDTH_IN_MAX <= 0) begin : gen_error_WIDTH_IN_MAX
            initial begin
                $error("DATA_WIDTH_IN_MAX must be > 0");
            end
        end

        if (WIDTH_OUT <= 0) begin : gen_error_WIDTH_OUT
            initial begin
                $error("DATA_WIDTH_OUT must be > 0");
            end
        end

        if (DIFFWIDTH < 0) begin : gen_error_DIFFWIDTH
            initial begin
                $error("WIDTH_OUT (%0d) cannot be larger than WIDTH_IN_MAX (%0d)",
                        WIDTH_OUT, WIDTH_IN_MAX);
            end
        end


        //=======================================================
        // If no bit difference, just pass through
        if (DIFFWIDTH == 0) begin : gen_pass_throught
            always_ff @(posedge clk) begin
                if (ena) begin
                    dout <=din_t;
                end
            end
        end
        else begin : gen_rounding
            logic signed [WIDTH_OUT-1:0]   d_rounded;
            logic signed [WIDTH_OUT-1:0]   d_trunc;
            logic                          round_up;
            logic signed [WIDTH_OUT:0]     d_temp; // one extra bit for rounding carry

            always_comb begin
                // Step 1: truncate to target width
                d_trunc =din_t[WIDTH_IN_MAX-1:DIFFWIDTH];

                // Step 2: unbiased rounding (round-half-to-even)
                round_up  = (din_t[DIFFWIDTH-1:0] > FRAC05) ||
                            ((din_t[DIFFWIDTH-1:0] == FRAC05) && d_trunc[0]);

                // 3. Apply rounding depending on mode
                if (IS_SIGNED) begin : gen_signed_rounding
                    // Signed rounding
                    d_temp = {d_trunc[WIDTH_OUT-1], d_trunc} +
                            (din_t[WIDTH_IN_MAX-1] ? -round_up : round_up);
                end
                else begin : gen_unsigned_rounding
                    // Unsigned rounding
                    d_temp = {1'b0, d_trunc} + round_up;
                end


                // Step 4: saturation check
                if (IS_SIGNED) begin : gen_signed_saturation
                    // Signed saturation
                    if (d_temp[WIDTH_OUT] != d_temp[WIDTH_OUT-1]) begin
                        // overflow happened
                        d_rounded =din_t[WIDTH_IN_MAX-1] ? MINVALsigned : MAXVALsigned;
                    end else begin
                        // no overflow
                        d_rounded = d_temp[WIDTH_OUT-1:0];
                    end
                end
                else begin : gen_unsigned_saturation
                    // Unsigned saturation
                    if (d_temp[WIDTH_OUT])
                        d_rounded = MAXVALunsigned;
                    else
                        d_rounded = d_temp[WIDTH_OUT-1:0];
                end
            end


            always_ff @(posedge clk) begin
                if (ena) begin
                    dout <= d_rounded;
                end
            end
        end
    endgenerate


    // (Synthesizers usually ignore 'initial' blocks for logic generation)
    initial begin
        if (width_in > WIDTH_OUT)
            $error("Parameter width_in must be <= WIDTH_OUT");
    end

endmodule
